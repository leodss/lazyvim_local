Vim�UnDo� �vG?JO����a�!�*1Ȯ��+
��į	   X     covergroup cg_val;                             fi�f    _�                            ����                                                                                                                                                                                                                                                                                                                                                             fi�f     �         X        covergroup cg_val;      5��                         e                     5�_�                            ����                                                                                                                                                                                                                                                                                                                                                             fi�b     �         X        covergroup cg_val;    5��                         e                     5��